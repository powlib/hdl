`ifndef POWLIB_IP 
`define POWLIB_IP

`define POWLIB_OPW      1    // Operation Width
`define POWLIB_OP_WRITE 1'd0 // Write Operation
`define POWLIB_OP_READ  1'd1 // Read Operation

`define AXI_LENW        8
`define AXI_SIZEW       3
`define AXI_BURSTW      2
`define AXI_RESPW       2
`define AXI_INCRBT      2d1

`endif