`ifndef POWLIB_IP 
`define POWLIB_IP

`define POWLIB_OPW      1 // Operation Width
`define POWLIB_OP_WRITE 0 // Write Operation
`define POWLIB_OP_READ  1 // Read Operation

`endif